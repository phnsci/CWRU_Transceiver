module CWRU_Transceiver_RX(
	inout [35:0] GPIO_1;
	output [6:0] HEX0
	);

endmodule