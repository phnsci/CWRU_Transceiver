module LED_display(input clk, code, output [6:0] HEX0);

always @(posedge clk)
begin
//	if (code == 'b01000000)
//		
//	else if (code == 'b01010000)
//		
//	else if (code == 'b01010100)
//		
//	else if (code == 'b01010101)
		
end

endmodule