module CWRU_Transceiver_RX(
	
	);

endmodule