`timescale 1 ns / 100 ps

module CWRU_Transceiver_RX_tb();



endmodule